library verilog;
use verilog.vl_types.all;
entity Registrador_vlg_vec_tst is
end Registrador_vlg_vec_tst;
