library verilog;
use verilog.vl_types.all;
entity Questao3 is
    port(
        gray            : in     vl_logic_vector(3 downto 0);
        johnson         : out    vl_logic_vector(4 downto 0)
    );
end Questao3;
