library verilog;
use verilog.vl_types.all;
entity Questao1b_vlg_vec_tst is
end Questao1b_vlg_vec_tst;
