library verilog;
use verilog.vl_types.all;
entity Mux_vlg_vec_tst is
end Mux_vlg_vec_tst;
