library verilog;
use verilog.vl_types.all;
entity Maquinas_vlg_check_tst is
    port(
        M1              : in     vl_logic;
        M2              : in     vl_logic;
        M3              : in     vl_logic;
        M4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Maquinas_vlg_check_tst;
