library verilog;
use verilog.vl_types.all;
entity Mux_vlg_check_tst is
    port(
        T               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Mux_vlg_check_tst;
