library verilog;
use verilog.vl_types.all;
entity Decodificador_vlg_vec_tst is
end Decodificador_vlg_vec_tst;
