library verilog;
use verilog.vl_types.all;
entity Questao1b_vlg_check_tst is
    port(
        X               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Questao1b_vlg_check_tst;
