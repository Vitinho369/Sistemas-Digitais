library verilog;
use verilog.vl_types.all;
entity Questao1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        x               : out    vl_logic
    );
end Questao1;
