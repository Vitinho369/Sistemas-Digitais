library verilog;
use verilog.vl_types.all;
entity Maquinas_vlg_vec_tst is
end Maquinas_vlg_vec_tst;
