library verilog;
use verilog.vl_types.all;
entity Questao1b is
    port(
        X               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic
    );
end Questao1b;
