library verilog;
use verilog.vl_types.all;
entity DecoderBCD_vlg_vec_tst is
end DecoderBCD_vlg_vec_tst;
