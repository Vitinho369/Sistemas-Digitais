library verilog;
use verilog.vl_types.all;
entity Questao3_vlg_check_tst is
    port(
        johnson         : in     vl_logic_vector(4 downto 0);
        sampler_rx      : in     vl_logic
    );
end Questao3_vlg_check_tst;
