library verilog;
use verilog.vl_types.all;
entity Questao5_vlg_vec_tst is
end Questao5_vlg_vec_tst;
