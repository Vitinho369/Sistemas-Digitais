library verilog;
use verilog.vl_types.all;
entity Questao3_vlg_sample_tst is
    port(
        gray            : in     vl_logic_vector(3 downto 0);
        sampler_tx      : out    vl_logic
    );
end Questao3_vlg_sample_tst;
