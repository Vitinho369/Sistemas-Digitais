library verilog;
use verilog.vl_types.all;
entity Subtrator_vlg_check_tst is
    port(
        s               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Subtrator_vlg_check_tst;
