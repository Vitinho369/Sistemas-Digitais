library verilog;
use verilog.vl_types.all;
entity Questao3_vlg_vec_tst is
end Questao3_vlg_vec_tst;
