library verilog;
use verilog.vl_types.all;
entity Questao1_vlg_vec_tst is
end Questao1_vlg_vec_tst;
