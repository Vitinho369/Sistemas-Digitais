library verilog;
use verilog.vl_types.all;
entity SeteSegmentos_vlg_vec_tst is
end SeteSegmentos_vlg_vec_tst;
